test_entity_name
  # (
    .a(a),
    .b(b),
    .c(c),
    .d(d),
    .e(e),
    .f(f)
  )

  test_entity_name_dut (
    g(g),
    h(h),
    i(i)
  );
